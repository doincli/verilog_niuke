`timescale 1ns / 1ps

 module phase_top    #(parameter DW=16) //   this is the top module;
(               
clk,
rst_n,
S1_data_in,
S2_data_in,
S1_data_tvaild,
S2_data_tvaild,
S1_data_out,
S2_data_out,
Number_w,
phase
);
/*** input and output ports ***/
input wire clk ;
input wire rst_n ;
input wire [DW-1:0] S1_data_in ;
input wire S1_data_tvaild ;
input wire S2_data_tvaild ;
input wire [DW-1:0] S2_data_in ;
output wire [DW-1:0] S1_data_out ;
output wire [DW-1:0] S2_data_out ; 
output wire [8:0] Number_w; 
output wire [18:0] phase;


/**************** wire and reg declaration *******************/

/*********** FFT wire and reg ******************/
wire [31:0]  S1_data_FFT ;
wire S1_data_FFT_tvalid ;
wire [15:0] S1_data_FFT_Re ;  // fix16_15 
wire [15:0] S1_data_FFT_Im ; // fix16_15 

wire [31:0]  S2_data_FFT ;
wire S2_data_FFT_tvalid ; 
wire [15:0]  S2_data_FFT_Re ; // fix16_15 
wire [15:0]  S2_data_FFT_Im ; // fix16_15 

wire [8:0] S1_index ;
wire [8:0] S2_index ;

reg FFT_cnt_en_S ;

reg [9:0] FFT_cnt_S ;  //  �������� FFT����ֻ��ȡ 512����Ч���ݣ�һ�����ڲ�����Ϊ512������ӦFFT����512����


/****** ��ģֵ��� wire ang reg ********/
wire [31:0] S1_data_FFT_Re2;  
wire [31:0] S1_data_FFT_Im2; 
wire [31:0] S2_data_FFT_Re2; 
wire [31:0] S2_data_FFT_Im2; 

wire [32:0] S1_data_FFT_module ; 
wire [32:0] S2_data_FFT_module ; 

/****** compare wire and reg ******/
wire [32:0]  S1_data_FFT_module_max;
wire [32:0]  S2_data_FFT_module_max;

reg [9:0] Location_S1;
reg [32:0] S1_data_FFT_module_1;
reg [32:0] S1_data_FFT_module_2;
reg [9:0] Location_S2;
reg [32:0] S2_data_FFT_module_1;
reg [32:0] S2_data_FFT_module_2;

/*****  arctan wire and reg ********/
reg [9:0] FFT_cnt_S1_1 ;  //  �������� arctan ������λ�ṩ���� ��������
reg [9:0] FFT_cnt_S2_1 ; 
wire      arctan_S1_en  ;
wire      arctan_S2_en  ;
reg      arctan_S1_en_reg  ;
reg      arctan_S2_en_reg  ;

wire  [17:0] phase_S1;
wire        phase_S1_vaild;
wire  [17:0] phase_S2;
wire        phase_S2_vaild;

/***** Number wire and reg *******/
wire  [18:0]  phase_S2_S1 ;
wire [18:0]  phase_step;
wire phase_Number_vaild; 
wire [47:0]  phase_out_data ;  
wire [17:0] phase_Number ;  //  �������֣�
wire [17:0]  little_data ;   //  С�����֣�

wire [23:0] phase_step_1 ;
wire [33:0] step ;

/****** phase_correction wire and reg ******/
reg [8:0] Number;
reg [15:0] S1_data_out_reg_1 ;
reg [15:0] S1_data_out_reg_2 ;
reg [15:0] S2_data_out_reg ;

reg [2047:0] data_out_1 ;
reg [2047:0] data_out_2 ;
reg [2047:0] data_out_3 ;
reg [2047:0] data_out_4 ;

reg [18:0] phase_g ;


assign S1_data_FFT_Im = S1_data_FFT[31:16];
assign S1_data_FFT_Re = S1_data_FFT[15:0] ;

assign S2_data_FFT_Im = S2_data_FFT[31:16];
assign S2_data_FFT_Re = S2_data_FFT[15:0] ;

always@(posedge clk) begin   //  �������ɼ��������� FFT����ֻ��ȡ 128����Ч����
     if(!rst_n) 
	    FFT_cnt_S <= 10'b0 ;		
	 else if(FFT_cnt_S== 10'd512)
	    FFT_cnt_S <=10'd512;  
     else if(S1_data_FFT_tvalid == 1'b1)	
        FFT_cnt_S <= FFT_cnt_S +10'b1 ;	 
	 else 
	    FFT_cnt_S <= 10'b0 ;	
end  

always@(posedge clk) begin  //  ��������cordic ���ݵ���Ч��ֵ 
     if(!rst_n)
        FFT_cnt_en_S <= 1'b0 ;
     else if(FFT_cnt_S == 10'd511) //== 8'd128) 
        FFT_cnt_en_S <= 1'b0 ;
     else if(FFT_cnt_S == 10'd512)//== 8'd129)
        FFT_cnt_en_S <= 1'b0 ;
     else if(S1_data_FFT_tvalid == 1'b1)
        FFT_cnt_en_S <= 1'b1 ;
     else 
        FFT_cnt_en_S <= 1'b0 ;
end


/*********** module1:�������źŵ� FFT �ķ�ֵ ***************/
FFT UU1_S1 (
  .aclk(clk),                                                // input wire aclk
  .aresetn(rst_n),                                          // input wire aresetn
  .s_axis_config_tdata(8'b1),                  // input wire [7 : 0] s_axis_config_tdata
  .s_axis_config_tvalid(1),                // input wire s_axis_config_tvalid
  .s_axis_config_tready(),                // output wire s_axis_config_tready
  .s_axis_data_tdata({16'b0,S1_data_in}),                      // input wire [31 : 0] s_axis_data_tdata
  .s_axis_data_tvalid(S1_data_tvaild),                    // input wire s_axis_data_tvalid
  .s_axis_data_tready(),                    // output wire s_axis_data_tready
  .s_axis_data_tlast(1),                      // input wire s_axis_data_tlast
  .m_axis_data_tdata(S1_data_FFT),                      // output wire [31 : 0] m_axis_data_tdata
  .m_axis_data_tuser(S1_index),                      // output wire [23 : 0] m_axis_data_tuser
  .m_axis_data_tvalid(S1_data_FFT_tvalid),                    // output wire m_axis_data_tvalid
  .m_axis_data_tready(1),                    // input wire m_axis_data_tready
  .m_axis_data_tlast(),                      // output wire m_axis_data_tlast
  .m_axis_status_tdata(),                  // output wire [7 : 0] m_axis_status_tdata
  .m_axis_status_tvalid(),                // output wire m_axis_status_tvalid
  .m_axis_status_tready(1),                // input wire m_axis_status_tready
  .event_frame_started(),                  // output wire event_frame_started
  .event_tlast_unexpected(),            // output wire event_tlast_unexpected
  .event_tlast_missing(),                  // output wire event_tlast_missing
  .event_status_channel_halt(),      // output wire event_status_channel_halt
  .event_data_in_channel_halt(),    // output wire event_data_in_channel_halt
  .event_data_out_channel_halt()  // output wire event_data_out_channel_halt
);

FFT UU1_S2 (
  .aclk(clk),                                                // input wire aclk
  .aresetn(rst_n),                                          // input wire aresetn
  .s_axis_config_tdata(8'b1),                  // input wire [7 : 0] s_axis_config_tdata
  .s_axis_config_tvalid(1),                // input wire s_axis_config_tvalid
  .s_axis_config_tready(),                // output wire s_axis_config_tready
  .s_axis_data_tdata({16'b0,S2_data_in}),                      // input wire [31 : 0] s_axis_data_tdata
  .s_axis_data_tvalid(S2_data_tvaild),                    // input wire s_axis_data_tvalid
  .s_axis_data_tready(),                    // output wire s_axis_data_tready
  .s_axis_data_tlast(1),                      // input wire s_axis_data_tlast
  .m_axis_data_tdata(S2_data_FFT),                      // output wire [31 : 0] m_axis_data_tdata
  .m_axis_data_tuser(S2_index),                      // output wire [23 : 0] m_axis_data_tuser
  .m_axis_data_tvalid(S2_data_FFT_tvalid),                    // output wire m_axis_data_tvalid
  .m_axis_data_tready(1),                    // input wire m_axis_data_tready
  .m_axis_data_tlast(),                      // output wire m_axis_data_tlast
  .m_axis_status_tdata(),                  // output wire [7 : 0] m_axis_status_tdata
  .m_axis_status_tvalid(),                // output wire m_axis_status_tvalid
  .m_axis_status_tready(1),                // input wire m_axis_status_tready
  .event_frame_started(),                  // output wire event_frame_started
  .event_tlast_unexpected(),            // output wire event_tlast_unexpected
  .event_tlast_missing(),                  // output wire event_tlast_missing
  .event_status_channel_halt(),      // output wire event_status_channel_halt
  .event_data_in_channel_halt(),    // output wire event_data_in_channel_halt
  .event_data_out_channel_halt()  // output wire event_data_out_channel_halt
);


/*********** module2: ��FFT ʵ���鲿�� ��ֵ  ���ó˷�����**************/ 
assign S1_data_FFT_module = {{S1_data_FFT_Re2[31]},S1_data_FFT_Re2}+{{S1_data_FFT_Im2[31]},S1_data_FFT_Im2};
assign S2_data_FFT_module = {{S2_data_FFT_Re2[31]},S2_data_FFT_Re2}+{{S2_data_FFT_Im2[31]},S2_data_FFT_Im2};

multiplier UU2_S1_RE (
  .CLK(clk),  // input wire CLK                   //  �����źſ���Ҫ���е���
  .A(S1_data_FFT_Re),      // input wire [15 : 0] A
  .B(S1_data_FFT_Re),      // input wire [15 : 0] B
  .P(S1_data_FFT_Re2)      // output wire [31 : 0] P
);
multiplier UU2_S1_IM (
  .CLK(clk),  // input wire CLK
  .A(S1_data_FFT_Im),      // input wire [15 : 0] A
  .B(S1_data_FFT_Im),      // input wire [15 : 0] B
  .P(S1_data_FFT_Im2)      // output wire [31 : 0] P
);
multiplier UU2_S2_RE (
  .CLK(clk),  // input wire CLK
  .A(S2_data_FFT_Re),      // input wire [15 : 0] A
  .B(S2_data_FFT_Re),      // input wire [15 : 0] B
  .P(S2_data_FFT_Re2)      // output wire [31 : 0] P
);
multiplier UU2_S2_IM (
  .CLK(clk),  // input wire CLK
  .A(S2_data_FFT_Im),      // input wire [15 : 0] A
  .B(S2_data_FFT_Im),      // input wire [15 : 0] B
  .P(S2_data_FFT_Im2)      // output wire [31 : 0] P
);


/********** module3: �Ƚ����ģֵ����ȡ��Ӧ��λ�� compare and location ***************/


compare  UU3_S1
(
.clk(clk),  //input wire clk_128M
.rst_n(rst_n),     //input wire rst_n 
.data0(S1_data_FFT_module),     //input wire [32:0] data0 
.FFT_cnt(FFT_cnt_S),   //input wire [9:0] FFT_cnt 
.FFT_cnt_en(FFT_cnt_en_S),  //input wire FFT_cnt_en
.data_max(S1_data_FFT_module_max)    //output wire [32:0] data_max 
);
compare  UU3_S2
(
.clk(clk),  //input wire clk_128M
.rst_n(rst_n),     //input wire rst_n 
.data0(S2_data_FFT_module),     //input wire [32:0] data0 
.FFT_cnt(FFT_cnt_S),   //input wire [9:0] FFT_cnt 
.FFT_cnt_en(FFT_cnt_en_S),  //input wire FFT_cnt_en
.data_max(S2_data_FFT_module_max)    //output wire [32:0] data_max 
);

always@(posedge clk) begin
   S1_data_FFT_module_1 <= S1_data_FFT_module;
   S1_data_FFT_module_2 <= S1_data_FFT_module_1;
   
   S2_data_FFT_module_1 <= S2_data_FFT_module;
   S2_data_FFT_module_2 <= S2_data_FFT_module_1;
end 

always@(posedge clk) begin
    if(!rst_n) 
	    Location_S1 <= 10'b0;
	else if(Location_S1) 
	    Location_S1 <= Location_S1;   
    else if(S1_data_FFT_module_max == 33'b0)  // Ϊ�˷�ֹ data_max ����Ϊ��󻹼������бȽ�
	    Location_S1 <= 10'b0;
    else if(S1_data_FFT_module_max == S1_data_FFT_module_2)
	    Location_S1 <= FFT_cnt_S - 10'd3;
    else 
        Location_S1 <= 10'b0;	   
end

always@(posedge clk) begin
    if(!rst_n) 
	    Location_S2 <= 10'b0;
	else if(Location_S2) 
        Location_S2 <= Location_S2;       
	else if(S2_data_FFT_module_max == 33'b0) // Ϊ�˷�ֹ data_max ����Ϊ��󻹼������бȽ�
        Location_S2 <= 10'b0;	
    else if(S2_data_FFT_module_max == S2_data_FFT_module_2)
	    Location_S2 <= FFT_cnt_S - 10'd3;
    else 
        Location_S2 <= 10'b0;	
end

/********** module3: ��S1��S2 ��λ�� arctan  **************/
assign arctan_S1_en = arctan_S1_en_reg ;
assign arctan_S2_en = arctan_S2_en_reg ;

always@(posedge clk) begin
    if(!rst_n) 
	    FFT_cnt_S1_1 <= 10'b0;
	else if(FFT_cnt_S1_1==10'd512) 
        FFT_cnt_S1_1 <= 10'd512;           
	else if(FFT_cnt_S==10'd510)
        FFT_cnt_S1_1 <= 10'b0; 
    else if(FFT_cnt_S==10'd512||FFT_cnt_S==10'd511) 
        FFT_cnt_S1_1 <= FFT_cnt_S1_1+10'b1;                
    else 
        FFT_cnt_S1_1 <= 10'b0;	
end

always@(posedge clk) begin
    if(!rst_n) 
	    FFT_cnt_S2_1 <= 10'b0;
	else if(FFT_cnt_S2_1==10'd512) 
        FFT_cnt_S2_1 <= 10'd512;           
	else if(FFT_cnt_S==10'd510)
        FFT_cnt_S2_1 <= 10'b0; 
    else if(FFT_cnt_S==10'd512||FFT_cnt_S==10'd511) 
        FFT_cnt_S2_1 <= FFT_cnt_S2_1+10'b1;                 
    else 
        FFT_cnt_S2_1 <= 10'b0;	
end

always@(posedge clk) begin
   if(!rst_n) 
      arctan_S1_en_reg <= 1'b0;
   else if((FFT_cnt_S1_1 == Location_S1) && Location_S1 )
      arctan_S1_en_reg <= 1'b1;
   else 
      arctan_S1_en_reg <= 1'b0;  
end

always@(posedge clk) begin
   if(!rst_n) 
      arctan_S2_en_reg <= 1'b0;
   else if((FFT_cnt_S2_1 == Location_S2) && Location_S2)
      arctan_S2_en_reg <= 1'b1;
   else 
      arctan_S2_en_reg <= 1'b0;  
end

arctan  UU4_S1(
  .aclk(clk),                                        // input wire aclk
  .s_axis_cartesian_tvalid(arctan_S1_en),  // input wire s_axis_cartesian_tvalid
  .s_axis_cartesian_tdata({{8{S1_data_FFT_Im[15]}},S1_data_FFT_Im,{8{S1_data_FFT_Re[15]}},S1_data_FFT_Re}), // input wire [47 : 0] s_axis_cartesian_tdata     
  .m_axis_dout_tvalid(phase_S1_vaild),            // output wire m_axis_dout_tvalid
  .m_axis_dout_tdata(phase_S1)              // output wire [23 : 0] m_axis_dout_tdata
);

arctan  UU4_S2(
  .aclk(clk),                                        // input wire aclk
  .s_axis_cartesian_tvalid(arctan_S2_en),  // input wire s_axis_cartesian_tvalid
  .s_axis_cartesian_tdata({{8{S2_data_FFT_Im[15]}},S2_data_FFT_Im,{8{S2_data_FFT_Re[15]}},S2_data_FFT_Re}), //  // input wire [47 : 0] s_axis_cartesian_tdata     
  .m_axis_dout_tvalid(phase_S2_vaild),            // output wire m_axis_dout_tvalid
  .m_axis_dout_tdata(phase_S2)              // output wire [23 : 0] m_axis_dout_tdata
);



/************* module4: ����λ�������Ҫ�Ĳ������� ***************/
assign  phase_S2_S1 = {phase_S2[17],phase_S2} - {phase_S1[17],phase_S1} ;  // fix 19_15

//assign  phase_step = 17'b00000000011001001;   fix17_14
assign  phase_step_1 = 24'b000000000011001001000011; // fix24_20

mult_gen_0 UU5_1 (     //  �������г���������Ƶ�ʵĵ���
  .CLK(clk),  // input wire CLK
  .A(phase_step_1),      // input wire [23 : 0] A
  .B(Location_S2),      // input wire [9 : 0] B
  .P(step)      // output wire [33 : 0] P
);
assign phase_step = step[23:5] ;

/*****************
������չ�� phase_step ��λ���� phase_step ��չ�� �˷����޵Ŀ�ȣ�
�ٶ���һ�� 17 bit λ������ݣ�
******************/

assign  phase_Number = phase_out_data[41:24];
assign  little_data  = phase_out_data[17:0];
phase_number UU5 (
  .aclk(clk),                                      // input wire aclk
  .s_axis_divisor_tvalid(1'b1),    // input wire s_axis_divisor_tvalid
  .s_axis_divisor_tdata({5'b0,phase_step}),      // input wire [23 : 0] s_axis_divisor_tdata
  .s_axis_dividend_tvalid(phase_S2_vaild),  // input wire s_axis_dividend_tvalid
  .s_axis_dividend_tdata({{5{phase_S2_S1[18]}},phase_S2_S1}),    // input wire [23 : 0] s_axis_dividend_tdata
  .m_axis_dout_tvalid(phase_Number_vaild),          // output wire m_axis_dout_tvalid
  .m_axis_dout_tdata(phase_out_data)            // output wire [47 : 0] m_axis_dout_tdata
);

assign phase = phase_g ;
always@(posedge clk) begin     //  ����λ����Ч����ס�������
   if(!rst_n) begin
      phase_g <= 19'b0 ;
   end
   else if(phase_S2_vaild) begin
      phase_g <= phase_S2_S1;
   end
   else begin
      phase_g <= phase_g ;
   end
end

/**************  module5: ͨ������������λ��������������λ���� *********************/

always@(posedge clk) begin    //ʹ�����ȡ��ֵ�����ֺ㶨��
   if(phase_Number_vaild)
   //if(phase_Number_vaild_1)
       Number <= phase_Number ;  
   else if(Number) 
       Number <= Number ;  //  �Ѳ����λ������������
   else 
       Number <= 9'b0 ;
end

assign S1_data_out = S1_data_out_reg_2 ; 
always@(posedge clk) begin  
   S1_data_out_reg_1 <= S1_data_in ;
   S1_data_out_reg_2 <= S1_data_out_reg_1 ;
end

always@(posedge clk) begin     // ͨ�������λ�������ʵ����ʱ������
   if(!rst_n) begin
      data_out_1 <=  2048'b0 ;
      data_out_2 <=  2048'b0 ;
      data_out_3 <=  2048'b0 ;
      data_out_4 <=  2048'b0 ;
   end
   else begin
       data_out_1 <=  {data_out_1[2031:0],S2_data_in} ;
       data_out_2 <=  {data_out_2[2031:0],data_out_1[2047:2032]} ;
       data_out_3 <=  {data_out_3[2031:0],data_out_2[2047:2032]} ;
       data_out_4 <=  {data_out_4[2031:0],data_out_3[2047:2032]} ;
    end       
end


assign S2_data_out = S2_data_out_reg ;
always@(posedge clk)  begin 
   case(Number)
   9'd0: begin S2_data_out_reg <= data_out_1[15:0]; end
   9'd1: begin S2_data_out_reg <= data_out_1[31:16]; end
   9'd2: begin S2_data_out_reg <= data_out_1[47:32]; end
   9'd3: begin S2_data_out_reg <= data_out_1[63:48]; end
   9'd4: begin S2_data_out_reg <= data_out_1[79:64]; end
   9'd5: begin S2_data_out_reg <= data_out_1[95:80]; end
   9'd6: begin S2_data_out_reg <= data_out_1[111:96]; end
   9'd7: begin S2_data_out_reg <= data_out_1[127:112]; end
   9'd8: begin S2_data_out_reg <= data_out_1[143:128]; end
   9'd9: begin S2_data_out_reg <= data_out_1[159:144]; end
   9'd10: begin S2_data_out_reg <= data_out_1[175:160]; end
   9'd11: begin S2_data_out_reg <= data_out_1[191:176]; end
   9'd12: begin S2_data_out_reg <= data_out_1[207:192]; end
   9'd13: begin S2_data_out_reg <= data_out_1[223:208]; end
   9'd14: begin S2_data_out_reg <= data_out_1[239:224]; end
   9'd15: begin S2_data_out_reg <= data_out_1[255:240]; end
   9'd16: begin S2_data_out_reg <= data_out_1[271:256]; end
   9'd17: begin S2_data_out_reg <= data_out_1[287:272]; end
   9'd18: begin S2_data_out_reg <= data_out_1[303:288]; end
   9'd19: begin S2_data_out_reg <= data_out_1[319:304]; end
   9'd20: begin S2_data_out_reg <= data_out_1[335:320]; end
   9'd21: begin S2_data_out_reg <= data_out_1[351:336]; end
   9'd22: begin S2_data_out_reg <= data_out_1[367:352]; end
   9'd23: begin S2_data_out_reg <= data_out_1[383:368]; end
   9'd24: begin S2_data_out_reg <= data_out_1[399:384]; end
   9'd25: begin S2_data_out_reg <= data_out_1[415:400]; end
   9'd26: begin S2_data_out_reg <= data_out_1[431:416]; end
   9'd27: begin S2_data_out_reg <= data_out_1[447:432]; end
   9'd28: begin S2_data_out_reg <= data_out_1[463:448]; end
   9'd29: begin S2_data_out_reg <= data_out_1[479:464]; end
   9'd30: begin S2_data_out_reg <= data_out_1[495:480]; end
   9'd31: begin S2_data_out_reg <= data_out_1[511:496]; end
   9'd32: begin S2_data_out_reg <= data_out_1[527:512]; end
   9'd33: begin S2_data_out_reg <= data_out_1[543:528]; end
   9'd34: begin S2_data_out_reg <= data_out_1[559:544]; end
   9'd35: begin S2_data_out_reg <= data_out_1[575:560]; end
   9'd36: begin S2_data_out_reg <= data_out_1[591:576]; end
   9'd37: begin S2_data_out_reg <= data_out_1[607:592]; end
   9'd38: begin S2_data_out_reg <= data_out_1[623:608]; end
   9'd39: begin S2_data_out_reg <= data_out_1[639:624]; end
   9'd40: begin S2_data_out_reg <= data_out_1[655:640]; end
   9'd41: begin S2_data_out_reg <= data_out_1[671:656]; end
   9'd42: begin S2_data_out_reg <= data_out_1[687:672]; end
   9'd43: begin S2_data_out_reg <= data_out_1[703:688]; end
   9'd44: begin S2_data_out_reg <= data_out_1[719:704]; end
   9'd45: begin S2_data_out_reg <= data_out_1[735:720]; end
   9'd46: begin S2_data_out_reg <= data_out_1[751:736]; end
   9'd47: begin S2_data_out_reg <= data_out_1[767:752]; end
   9'd48: begin S2_data_out_reg <= data_out_1[783:768]; end
   9'd49: begin S2_data_out_reg <= data_out_1[799:784]; end
   9'd50: begin S2_data_out_reg <= data_out_1[815:800]; end
   9'd51: begin S2_data_out_reg <= data_out_1[831:816]; end
   9'd52: begin S2_data_out_reg <= data_out_1[847:832]; end
   9'd53: begin S2_data_out_reg <= data_out_1[863:848]; end
   9'd54: begin S2_data_out_reg <= data_out_1[879:864]; end
   9'd55: begin S2_data_out_reg <= data_out_1[895:880]; end
   9'd56: begin S2_data_out_reg <= data_out_1[911:896]; end
   9'd57: begin S2_data_out_reg <= data_out_1[927:912]; end
   9'd58: begin S2_data_out_reg <= data_out_1[943:928]; end
   9'd59: begin S2_data_out_reg <= data_out_1[959:944]; end
   9'd60: begin S2_data_out_reg <= data_out_1[975:960]; end
   9'd61: begin S2_data_out_reg <= data_out_1[991:976]; end
   9'd62: begin S2_data_out_reg <= data_out_1[1007:992]; end
   9'd63: begin S2_data_out_reg <= data_out_1[1023:1008]; end
   9'd64: begin S2_data_out_reg <= data_out_1[1039:1024]; end
   9'd65: begin S2_data_out_reg <= data_out_1[1055:1040]; end
   9'd66: begin S2_data_out_reg <= data_out_1[1071:1056]; end
   9'd67: begin S2_data_out_reg <= data_out_1[1087:1072]; end
   9'd68: begin S2_data_out_reg <= data_out_1[1103:1088]; end
   9'd69: begin S2_data_out_reg <= data_out_1[1119:1104]; end
   9'd70: begin S2_data_out_reg <= data_out_1[1135:1120]; end
   9'd71: begin S2_data_out_reg <= data_out_1[1151:1136]; end
   9'd72: begin S2_data_out_reg <= data_out_1[1167:1152]; end
   9'd73: begin S2_data_out_reg <= data_out_1[1183:1168]; end
   9'd74: begin S2_data_out_reg <= data_out_1[1199:1184]; end
   9'd75: begin S2_data_out_reg <= data_out_1[1215:1200]; end
   9'd76: begin S2_data_out_reg <= data_out_1[1231:1216]; end
   9'd77: begin S2_data_out_reg <= data_out_1[1247:1232]; end
   9'd78: begin S2_data_out_reg <= data_out_1[1263:1248]; end
   9'd79: begin S2_data_out_reg <= data_out_1[1279:1264]; end
   9'd80: begin S2_data_out_reg <= data_out_1[1295:1280]; end
   9'd81: begin S2_data_out_reg <= data_out_1[1311:1296]; end
   9'd82: begin S2_data_out_reg <= data_out_1[1327:1312]; end
   9'd83: begin S2_data_out_reg <= data_out_1[1343:1328]; end
   9'd84: begin S2_data_out_reg <= data_out_1[1359:1344]; end
   9'd85: begin S2_data_out_reg <= data_out_1[1375:1360]; end
   9'd86: begin S2_data_out_reg <= data_out_1[1391:1376]; end
   9'd87: begin S2_data_out_reg <= data_out_1[1407:1392]; end
   9'd88: begin S2_data_out_reg <= data_out_1[1423:1408]; end
   9'd89: begin S2_data_out_reg <= data_out_1[1439:1424]; end
   9'd90: begin S2_data_out_reg <= data_out_1[1455:1440]; end
   9'd91: begin S2_data_out_reg <= data_out_1[1471:1456]; end
   9'd92: begin S2_data_out_reg <= data_out_1[1487:1472]; end
   9'd93: begin S2_data_out_reg <= data_out_1[1503:1488]; end
   9'd94: begin S2_data_out_reg <= data_out_1[1519:1504]; end
   9'd95: begin S2_data_out_reg <= data_out_1[1535:1520]; end
   9'd96: begin S2_data_out_reg <= data_out_1[1551:1536]; end
   9'd97: begin S2_data_out_reg <= data_out_1[1567:1552]; end
   9'd98: begin S2_data_out_reg <= data_out_1[1583:1568]; end
   9'd99: begin S2_data_out_reg <= data_out_1[1599:1584]; end
   9'd100: begin S2_data_out_reg <= data_out_1[1615:1600]; end
   9'd101: begin S2_data_out_reg <= data_out_1[1631:1616]; end
   9'd102: begin S2_data_out_reg <= data_out_1[1647:1632]; end
   9'd103: begin S2_data_out_reg <= data_out_1[1663:1648]; end
   9'd104: begin S2_data_out_reg <= data_out_1[1679:1664]; end
   9'd105: begin S2_data_out_reg <= data_out_1[1695:1680]; end
   9'd106: begin S2_data_out_reg <= data_out_1[1711:1696]; end
   9'd107: begin S2_data_out_reg <= data_out_1[1727:1712]; end
   9'd108: begin S2_data_out_reg <= data_out_1[1743:1728]; end
   9'd109: begin S2_data_out_reg <= data_out_1[1759:1744]; end
   9'd110: begin S2_data_out_reg <= data_out_1[1775:1760]; end
   9'd111: begin S2_data_out_reg <= data_out_1[1791:1776]; end
   9'd112: begin S2_data_out_reg <= data_out_1[1807:1792]; end
   9'd113: begin S2_data_out_reg <= data_out_1[1823:1808]; end
   9'd114: begin S2_data_out_reg <= data_out_1[1839:1824]; end
   9'd115: begin S2_data_out_reg <= data_out_1[1855:1840]; end
   9'd116: begin S2_data_out_reg <= data_out_1[1871:1856]; end
   9'd117: begin S2_data_out_reg <= data_out_1[1887:1872]; end
   9'd118: begin S2_data_out_reg <= data_out_1[1903:1888]; end
   9'd119: begin S2_data_out_reg <= data_out_1[1919:1904]; end
   9'd120: begin S2_data_out_reg <= data_out_1[1935:1920]; end
   9'd121: begin S2_data_out_reg <= data_out_1[1951:1936]; end
   9'd122: begin S2_data_out_reg <= data_out_1[1967:1952]; end
   9'd123: begin S2_data_out_reg <= data_out_1[1983:1968]; end
   9'd124: begin S2_data_out_reg <= data_out_1[1999:1984]; end
   9'd125: begin S2_data_out_reg <= data_out_1[2015:2000]; end
   9'd126: begin S2_data_out_reg <= data_out_1[2031:2016]; end
   9'd127: begin S2_data_out_reg <= data_out_1[2047:2032]; end
   9'd128: begin S2_data_out_reg <= data_out_2[15:0]; end
   9'd129: begin S2_data_out_reg <= data_out_2[31:16]; end
   9'd130: begin S2_data_out_reg <= data_out_2[47:32]; end
   9'd131: begin S2_data_out_reg <= data_out_2[63:48]; end
   9'd132: begin S2_data_out_reg <= data_out_2[79:64]; end
   9'd133: begin S2_data_out_reg <= data_out_2[95:80]; end
   9'd134: begin S2_data_out_reg <= data_out_2[111:96]; end
   9'd135: begin S2_data_out_reg <= data_out_2[127:112]; end
   9'd136: begin S2_data_out_reg <= data_out_2[143:128]; end
   9'd137: begin S2_data_out_reg <= data_out_2[159:144]; end
   9'd138: begin S2_data_out_reg <= data_out_2[175:160]; end
   9'd139: begin S2_data_out_reg <= data_out_2[191:176]; end
   9'd140: begin S2_data_out_reg <= data_out_2[207:192]; end
   9'd141: begin S2_data_out_reg <= data_out_2[223:208]; end
   9'd142: begin S2_data_out_reg <= data_out_2[239:224]; end
   9'd143: begin S2_data_out_reg <= data_out_2[255:240]; end
   9'd144: begin S2_data_out_reg <= data_out_2[271:256]; end
   9'd145: begin S2_data_out_reg <= data_out_2[287:272]; end
   9'd146: begin S2_data_out_reg <= data_out_2[303:288]; end
   9'd147: begin S2_data_out_reg <= data_out_2[319:304]; end
   9'd148: begin S2_data_out_reg <= data_out_2[335:320]; end
   9'd149: begin S2_data_out_reg <= data_out_2[351:336]; end
   9'd150: begin S2_data_out_reg <= data_out_2[367:352]; end
   9'd151: begin S2_data_out_reg <= data_out_2[383:368]; end
   9'd152: begin S2_data_out_reg <= data_out_2[399:384]; end
   9'd153: begin S2_data_out_reg <= data_out_2[415:400]; end
   9'd154: begin S2_data_out_reg <= data_out_2[431:416]; end
   9'd155: begin S2_data_out_reg <= data_out_2[447:432]; end
   9'd156: begin S2_data_out_reg <= data_out_2[463:448]; end
   9'd157: begin S2_data_out_reg <= data_out_2[479:464]; end
   9'd158: begin S2_data_out_reg <= data_out_2[495:480]; end
   9'd159: begin S2_data_out_reg <= data_out_2[511:496]; end
   9'd160: begin S2_data_out_reg <= data_out_2[527:512]; end
   9'd161: begin S2_data_out_reg <= data_out_2[543:528]; end
   9'd162: begin S2_data_out_reg <= data_out_2[559:544]; end
   9'd163: begin S2_data_out_reg <= data_out_2[575:560]; end
   9'd164: begin S2_data_out_reg <= data_out_2[591:576]; end
   9'd165: begin S2_data_out_reg <= data_out_2[607:592]; end
   9'd166: begin S2_data_out_reg <= data_out_2[623:608]; end
   9'd167: begin S2_data_out_reg <= data_out_2[639:624]; end
   9'd168: begin S2_data_out_reg <= data_out_2[655:640]; end
   9'd169: begin S2_data_out_reg <= data_out_2[671:656]; end
   9'd170: begin S2_data_out_reg <= data_out_2[687:672]; end
   9'd171: begin S2_data_out_reg <= data_out_2[703:688]; end
   9'd172: begin S2_data_out_reg <= data_out_2[719:704]; end
   9'd173: begin S2_data_out_reg <= data_out_2[735:720]; end
   9'd174: begin S2_data_out_reg <= data_out_2[751:736]; end
   9'd175: begin S2_data_out_reg <= data_out_2[767:752]; end
   9'd176: begin S2_data_out_reg <= data_out_2[783:768]; end
   9'd177: begin S2_data_out_reg <= data_out_2[799:784]; end
   9'd178: begin S2_data_out_reg <= data_out_2[815:800]; end
   9'd179: begin S2_data_out_reg <= data_out_2[831:816]; end
   9'd180: begin S2_data_out_reg <= data_out_2[847:832]; end
   9'd181: begin S2_data_out_reg <= data_out_2[863:848]; end
   9'd182: begin S2_data_out_reg <= data_out_2[879:864]; end
   9'd183: begin S2_data_out_reg <= data_out_2[895:880]; end
   9'd184: begin S2_data_out_reg <= data_out_2[911:896]; end
   9'd185: begin S2_data_out_reg <= data_out_2[927:912]; end
   9'd186: begin S2_data_out_reg <= data_out_2[943:928]; end
   9'd187: begin S2_data_out_reg <= data_out_2[959:944]; end
   9'd188: begin S2_data_out_reg <= data_out_2[975:960]; end
   9'd189: begin S2_data_out_reg <= data_out_2[991:976]; end
   9'd190: begin S2_data_out_reg <= data_out_2[1007:992]; end
   9'd191: begin S2_data_out_reg <= data_out_2[1023:1008]; end
   9'd192: begin S2_data_out_reg <= data_out_2[1039:1024]; end
   9'd193: begin S2_data_out_reg <= data_out_2[1055:1040]; end
   9'd194: begin S2_data_out_reg <= data_out_2[1071:1056]; end
   9'd195: begin S2_data_out_reg <= data_out_2[1087:1072]; end
   9'd196: begin S2_data_out_reg <= data_out_2[1103:1088]; end
   9'd197: begin S2_data_out_reg <= data_out_2[1119:1104]; end
   9'd198: begin S2_data_out_reg <= data_out_2[1135:1120]; end
   9'd199: begin S2_data_out_reg <= data_out_2[1151:1136]; end
   9'd200: begin S2_data_out_reg <= data_out_2[1167:1152]; end
   9'd201: begin S2_data_out_reg <= data_out_2[1183:1168]; end
   9'd202: begin S2_data_out_reg <= data_out_2[1199:1184]; end
   9'd203: begin S2_data_out_reg <= data_out_2[1215:1200]; end
   9'd204: begin S2_data_out_reg <= data_out_2[1231:1216]; end
   9'd205: begin S2_data_out_reg <= data_out_2[1247:1232]; end
   9'd206: begin S2_data_out_reg <= data_out_2[1263:1248]; end
   9'd207: begin S2_data_out_reg <= data_out_2[1279:1264]; end
   9'd208: begin S2_data_out_reg <= data_out_2[1295:1280]; end
   9'd209: begin S2_data_out_reg <= data_out_2[1311:1296]; end
   9'd210: begin S2_data_out_reg <= data_out_2[1327:1312]; end
   9'd211: begin S2_data_out_reg <= data_out_2[1343:1328]; end
   9'd212: begin S2_data_out_reg <= data_out_2[1359:1344]; end
   9'd213: begin S2_data_out_reg <= data_out_2[1375:1360]; end
   9'd214: begin S2_data_out_reg <= data_out_2[1391:1376]; end
   9'd215: begin S2_data_out_reg <= data_out_2[1407:1392]; end
   9'd216: begin S2_data_out_reg <= data_out_2[1423:1408]; end
   9'd217: begin S2_data_out_reg <= data_out_2[1439:1424]; end
   9'd218: begin S2_data_out_reg <= data_out_2[1455:1440]; end
   9'd219: begin S2_data_out_reg <= data_out_2[1471:1456]; end
   9'd220: begin S2_data_out_reg <= data_out_2[1487:1472]; end
   9'd221: begin S2_data_out_reg <= data_out_2[1503:1488]; end
   9'd222: begin S2_data_out_reg <= data_out_2[1519:1504]; end
   9'd223: begin S2_data_out_reg <= data_out_2[1535:1520]; end
   9'd224: begin S2_data_out_reg <= data_out_2[1551:1536]; end
   9'd225: begin S2_data_out_reg <= data_out_2[1567:1552]; end
   9'd226: begin S2_data_out_reg <= data_out_2[1583:1568]; end
   9'd227: begin S2_data_out_reg <= data_out_2[1599:1584]; end
   9'd228: begin S2_data_out_reg <= data_out_2[1615:1600]; end
   9'd229: begin S2_data_out_reg <= data_out_2[1631:1616]; end
   9'd230: begin S2_data_out_reg <= data_out_2[1647:1632]; end
   9'd231: begin S2_data_out_reg <= data_out_2[1663:1648]; end
   9'd232: begin S2_data_out_reg <= data_out_2[1679:1664]; end
   9'd233: begin S2_data_out_reg <= data_out_2[1695:1680]; end
   9'd234: begin S2_data_out_reg <= data_out_2[1711:1696]; end
   9'd235: begin S2_data_out_reg <= data_out_2[1727:1712]; end
   9'd236: begin S2_data_out_reg <= data_out_2[1743:1728]; end
   9'd237: begin S2_data_out_reg <= data_out_2[1759:1744]; end
   9'd238: begin S2_data_out_reg <= data_out_2[1775:1760]; end
   9'd239: begin S2_data_out_reg <= data_out_2[1791:1776]; end
   9'd240: begin S2_data_out_reg <= data_out_2[1807:1792]; end
   9'd241: begin S2_data_out_reg <= data_out_2[1823:1808]; end
   9'd242: begin S2_data_out_reg <= data_out_2[1839:1824]; end
   9'd243: begin S2_data_out_reg <= data_out_2[1855:1840]; end
   9'd244: begin S2_data_out_reg <= data_out_2[1871:1856]; end
   9'd245: begin S2_data_out_reg <= data_out_2[1887:1872]; end
   9'd246: begin S2_data_out_reg <= data_out_2[1903:1888]; end
   9'd247: begin S2_data_out_reg <= data_out_2[1919:1904]; end
   9'd248: begin S2_data_out_reg <= data_out_2[1935:1920]; end
   9'd249: begin S2_data_out_reg <= data_out_2[1951:1936]; end
   9'd250: begin S2_data_out_reg <= data_out_2[1967:1952]; end
   9'd251: begin S2_data_out_reg <= data_out_2[1983:1968]; end
   9'd252: begin S2_data_out_reg <= data_out_2[1999:1984]; end
   9'd253: begin S2_data_out_reg <= data_out_2[2015:2000]; end
   9'd254: begin S2_data_out_reg <= data_out_2[2031:2016]; end
   9'd255: begin S2_data_out_reg <= data_out_2[2047:2032]; end
   9'd256: begin S2_data_out_reg <= data_out_3[15:0]; end
   9'd257: begin S2_data_out_reg <= data_out_3[31:16]; end
   9'd258: begin S2_data_out_reg <= data_out_3[47:32]; end
   9'd259: begin S2_data_out_reg <= data_out_3[63:48]; end
   9'd260: begin S2_data_out_reg <= data_out_3[79:64]; end
   9'd261: begin S2_data_out_reg <= data_out_3[95:80]; end
   9'd262: begin S2_data_out_reg <= data_out_3[111:96]; end
   9'd263: begin S2_data_out_reg <= data_out_3[127:112]; end
   9'd264: begin S2_data_out_reg <= data_out_3[143:128]; end
   9'd265: begin S2_data_out_reg <= data_out_3[159:144]; end
   9'd266: begin S2_data_out_reg <= data_out_3[175:160]; end
   9'd267: begin S2_data_out_reg <= data_out_3[191:176]; end
   9'd268: begin S2_data_out_reg <= data_out_3[207:192]; end
   9'd269: begin S2_data_out_reg <= data_out_3[223:208]; end
   9'd270: begin S2_data_out_reg <= data_out_3[239:224]; end
   9'd271: begin S2_data_out_reg <= data_out_3[255:240]; end
   9'd272: begin S2_data_out_reg <= data_out_3[271:256]; end
   9'd273: begin S2_data_out_reg <= data_out_3[287:272]; end
   9'd274: begin S2_data_out_reg <= data_out_3[303:288]; end
   9'd275: begin S2_data_out_reg <= data_out_3[319:304]; end
   9'd276: begin S2_data_out_reg <= data_out_3[335:320]; end
   9'd277: begin S2_data_out_reg <= data_out_3[351:336]; end
   9'd278: begin S2_data_out_reg <= data_out_3[367:352]; end
   9'd279: begin S2_data_out_reg <= data_out_3[383:368]; end
   9'd280: begin S2_data_out_reg <= data_out_3[399:384]; end
   9'd281: begin S2_data_out_reg <= data_out_3[415:400]; end
   9'd282: begin S2_data_out_reg <= data_out_3[431:416]; end
   9'd283: begin S2_data_out_reg <= data_out_3[447:432]; end
   9'd284: begin S2_data_out_reg <= data_out_3[463:448]; end
   9'd285: begin S2_data_out_reg <= data_out_3[479:464]; end
   9'd286: begin S2_data_out_reg <= data_out_3[495:480]; end
   9'd287: begin S2_data_out_reg <= data_out_3[511:496]; end
   9'd288: begin S2_data_out_reg <= data_out_3[527:512]; end
   9'd289: begin S2_data_out_reg <= data_out_3[543:528]; end
   9'd290: begin S2_data_out_reg <= data_out_3[559:544]; end
   9'd291: begin S2_data_out_reg <= data_out_3[575:560]; end
   9'd292: begin S2_data_out_reg <= data_out_3[591:576]; end
   9'd293: begin S2_data_out_reg <= data_out_3[607:592]; end
   9'd294: begin S2_data_out_reg <= data_out_3[623:608]; end
   9'd295: begin S2_data_out_reg <= data_out_3[639:624]; end
   9'd296: begin S2_data_out_reg <= data_out_3[655:640]; end
   9'd297: begin S2_data_out_reg <= data_out_3[671:656]; end
   9'd298: begin S2_data_out_reg <= data_out_3[687:672]; end
   9'd299: begin S2_data_out_reg <= data_out_3[703:688]; end
   9'd300: begin S2_data_out_reg <= data_out_3[719:704]; end
   9'd301: begin S2_data_out_reg <= data_out_3[735:720]; end
   9'd302: begin S2_data_out_reg <= data_out_3[751:736]; end
   9'd303: begin S2_data_out_reg <= data_out_3[767:752]; end
   9'd304: begin S2_data_out_reg <= data_out_3[783:768]; end
   9'd305: begin S2_data_out_reg <= data_out_3[799:784]; end
   9'd306: begin S2_data_out_reg <= data_out_3[815:800]; end
   9'd307: begin S2_data_out_reg <= data_out_3[831:816]; end
   9'd308: begin S2_data_out_reg <= data_out_3[847:832]; end
   9'd309: begin S2_data_out_reg <= data_out_3[863:848]; end
   9'd310: begin S2_data_out_reg <= data_out_3[879:864]; end
   9'd311: begin S2_data_out_reg <= data_out_3[895:880]; end
   9'd312: begin S2_data_out_reg <= data_out_3[911:896]; end
   9'd313: begin S2_data_out_reg <= data_out_3[927:912]; end
   9'd314: begin S2_data_out_reg <= data_out_3[943:928]; end
   9'd315: begin S2_data_out_reg <= data_out_3[959:944]; end
   9'd316: begin S2_data_out_reg <= data_out_3[975:960]; end
   9'd317: begin S2_data_out_reg <= data_out_3[991:976]; end
   9'd318: begin S2_data_out_reg <= data_out_3[1007:992]; end
   9'd319: begin S2_data_out_reg <= data_out_3[1023:1008]; end
   9'd320: begin S2_data_out_reg <= data_out_3[1039:1024]; end
   9'd321: begin S2_data_out_reg <= data_out_3[1055:1040]; end
   9'd322: begin S2_data_out_reg <= data_out_3[1071:1056]; end
   9'd323: begin S2_data_out_reg <= data_out_3[1087:1072]; end
   9'd324: begin S2_data_out_reg <= data_out_3[1103:1088]; end
   9'd325: begin S2_data_out_reg <= data_out_3[1119:1104]; end
   9'd326: begin S2_data_out_reg <= data_out_3[1135:1120]; end
   9'd327: begin S2_data_out_reg <= data_out_3[1151:1136]; end
   9'd328: begin S2_data_out_reg <= data_out_3[1167:1152]; end
   9'd329: begin S2_data_out_reg <= data_out_3[1183:1168]; end
   9'd330: begin S2_data_out_reg <= data_out_3[1199:1184]; end
   9'd331: begin S2_data_out_reg <= data_out_3[1215:1200]; end
   9'd332: begin S2_data_out_reg <= data_out_3[1231:1216]; end
   9'd333: begin S2_data_out_reg <= data_out_3[1247:1232]; end
   9'd334: begin S2_data_out_reg <= data_out_3[1263:1248]; end
   9'd335: begin S2_data_out_reg <= data_out_3[1279:1264]; end
   9'd336: begin S2_data_out_reg <= data_out_3[1295:1280]; end
   9'd337: begin S2_data_out_reg <= data_out_3[1311:1296]; end
   9'd338: begin S2_data_out_reg <= data_out_3[1327:1312]; end
   9'd339: begin S2_data_out_reg <= data_out_3[1343:1328]; end
   9'd340: begin S2_data_out_reg <= data_out_3[1359:1344]; end
   9'd341: begin S2_data_out_reg <= data_out_3[1375:1360]; end
   9'd342: begin S2_data_out_reg <= data_out_3[1391:1376]; end
   9'd343: begin S2_data_out_reg <= data_out_3[1407:1392]; end
   9'd344: begin S2_data_out_reg <= data_out_3[1423:1408]; end
   9'd345: begin S2_data_out_reg <= data_out_3[1439:1424]; end
   9'd346: begin S2_data_out_reg <= data_out_3[1455:1440]; end
   9'd347: begin S2_data_out_reg <= data_out_3[1471:1456]; end
   9'd348: begin S2_data_out_reg <= data_out_3[1487:1472]; end
   9'd349: begin S2_data_out_reg <= data_out_3[1503:1488]; end
   9'd350: begin S2_data_out_reg <= data_out_3[1519:1504]; end
   9'd351: begin S2_data_out_reg <= data_out_3[1535:1520]; end
   9'd352: begin S2_data_out_reg <= data_out_3[1551:1536]; end
   9'd353: begin S2_data_out_reg <= data_out_3[1567:1552]; end
   9'd354: begin S2_data_out_reg <= data_out_3[1583:1568]; end
   9'd355: begin S2_data_out_reg <= data_out_3[1599:1584]; end
   9'd356: begin S2_data_out_reg <= data_out_3[1615:1600]; end
   9'd357: begin S2_data_out_reg <= data_out_3[1631:1616]; end
   9'd358: begin S2_data_out_reg <= data_out_3[1647:1632]; end
   9'd359: begin S2_data_out_reg <= data_out_3[1663:1648]; end
   9'd360: begin S2_data_out_reg <= data_out_3[1679:1664]; end
   9'd361: begin S2_data_out_reg <= data_out_3[1695:1680]; end
   9'd362: begin S2_data_out_reg <= data_out_3[1711:1696]; end
   9'd363: begin S2_data_out_reg <= data_out_3[1727:1712]; end
   9'd364: begin S2_data_out_reg <= data_out_3[1743:1728]; end
   9'd365: begin S2_data_out_reg <= data_out_3[1759:1744]; end
   9'd366: begin S2_data_out_reg <= data_out_3[1775:1760]; end
   9'd367: begin S2_data_out_reg <= data_out_3[1791:1776]; end
   9'd368: begin S2_data_out_reg <= data_out_3[1807:1792]; end
   9'd369: begin S2_data_out_reg <= data_out_3[1823:1808]; end
   9'd370: begin S2_data_out_reg <= data_out_3[1839:1824]; end
   9'd371: begin S2_data_out_reg <= data_out_3[1855:1840]; end
   9'd372: begin S2_data_out_reg <= data_out_3[1871:1856]; end
   9'd373: begin S2_data_out_reg <= data_out_3[1887:1872]; end
   9'd374: begin S2_data_out_reg <= data_out_3[1903:1888]; end
   9'd375: begin S2_data_out_reg <= data_out_3[1919:1904]; end
   9'd376: begin S2_data_out_reg <= data_out_3[1935:1920]; end
   9'd377: begin S2_data_out_reg <= data_out_3[1951:1936]; end
   9'd378: begin S2_data_out_reg <= data_out_3[1967:1952]; end
   9'd379: begin S2_data_out_reg <= data_out_3[1983:1968]; end
   9'd380: begin S2_data_out_reg <= data_out_3[1999:1984]; end
   9'd381: begin S2_data_out_reg <= data_out_3[2015:2000]; end
   9'd382: begin S2_data_out_reg <= data_out_3[2031:2016]; end
   9'd383: begin S2_data_out_reg <= data_out_3[2047:2032]; end
   9'd384: begin S2_data_out_reg <= data_out_4[15:0]; end
   9'd385: begin S2_data_out_reg <= data_out_4[31:16]; end
   9'd386: begin S2_data_out_reg <= data_out_4[47:32]; end
   9'd387: begin S2_data_out_reg <= data_out_4[63:48]; end
   9'd388: begin S2_data_out_reg <= data_out_4[79:64]; end
   9'd389: begin S2_data_out_reg <= data_out_4[95:80]; end
   9'd390: begin S2_data_out_reg <= data_out_4[111:96]; end
   9'd391: begin S2_data_out_reg <= data_out_4[127:112]; end
   9'd392: begin S2_data_out_reg <= data_out_4[143:128]; end
   9'd393: begin S2_data_out_reg <= data_out_4[159:144]; end
   9'd394: begin S2_data_out_reg <= data_out_4[175:160]; end
   9'd395: begin S2_data_out_reg <= data_out_4[191:176]; end
   9'd396: begin S2_data_out_reg <= data_out_4[207:192]; end
   9'd397: begin S2_data_out_reg <= data_out_4[223:208]; end
   9'd398: begin S2_data_out_reg <= data_out_4[239:224]; end
   9'd399: begin S2_data_out_reg <= data_out_4[255:240]; end
   9'd400: begin S2_data_out_reg <= data_out_4[271:256]; end
   9'd401: begin S2_data_out_reg <= data_out_4[287:272]; end
   9'd402: begin S2_data_out_reg <= data_out_4[303:288]; end
   9'd403: begin S2_data_out_reg <= data_out_4[319:304]; end
   9'd404: begin S2_data_out_reg <= data_out_4[335:320]; end
   9'd405: begin S2_data_out_reg <= data_out_4[351:336]; end
   9'd406: begin S2_data_out_reg <= data_out_4[367:352]; end
   9'd407: begin S2_data_out_reg <= data_out_4[383:368]; end
   9'd408: begin S2_data_out_reg <= data_out_4[399:384]; end
   9'd409: begin S2_data_out_reg <= data_out_4[415:400]; end
   9'd410: begin S2_data_out_reg <= data_out_4[431:416]; end
   9'd411: begin S2_data_out_reg <= data_out_4[447:432]; end
   9'd412: begin S2_data_out_reg <= data_out_4[463:448]; end
   9'd413: begin S2_data_out_reg <= data_out_4[479:464]; end
   9'd414: begin S2_data_out_reg <= data_out_4[495:480]; end
   9'd415: begin S2_data_out_reg <= data_out_4[511:496]; end
   9'd416: begin S2_data_out_reg <= data_out_4[527:512]; end
   9'd417: begin S2_data_out_reg <= data_out_4[543:528]; end
   9'd418: begin S2_data_out_reg <= data_out_4[559:544]; end
   9'd419: begin S2_data_out_reg <= data_out_4[575:560]; end
   9'd420: begin S2_data_out_reg <= data_out_4[591:576]; end
   9'd421: begin S2_data_out_reg <= data_out_4[607:592]; end
   9'd422: begin S2_data_out_reg <= data_out_4[623:608]; end
   9'd423: begin S2_data_out_reg <= data_out_4[639:624]; end
   9'd424: begin S2_data_out_reg <= data_out_4[655:640]; end
   9'd425: begin S2_data_out_reg <= data_out_4[671:656]; end
   9'd426: begin S2_data_out_reg <= data_out_4[687:672]; end
   9'd427: begin S2_data_out_reg <= data_out_4[703:688]; end
   9'd428: begin S2_data_out_reg <= data_out_4[719:704]; end
   9'd429: begin S2_data_out_reg <= data_out_4[735:720]; end
   9'd430: begin S2_data_out_reg <= data_out_4[751:736]; end
   9'd431: begin S2_data_out_reg <= data_out_4[767:752]; end
   9'd432: begin S2_data_out_reg <= data_out_4[783:768]; end
   9'd433: begin S2_data_out_reg <= data_out_4[799:784]; end
   9'd434: begin S2_data_out_reg <= data_out_4[815:800]; end
   9'd435: begin S2_data_out_reg <= data_out_4[831:816]; end
   9'd436: begin S2_data_out_reg <= data_out_4[847:832]; end
   9'd437: begin S2_data_out_reg <= data_out_4[863:848]; end
   9'd438: begin S2_data_out_reg <= data_out_4[879:864]; end
   9'd439: begin S2_data_out_reg <= data_out_4[895:880]; end
   9'd440: begin S2_data_out_reg <= data_out_4[911:896]; end
   9'd441: begin S2_data_out_reg <= data_out_4[927:912]; end
   9'd442: begin S2_data_out_reg <= data_out_4[943:928]; end
   9'd443: begin S2_data_out_reg <= data_out_4[959:944]; end
   9'd444: begin S2_data_out_reg <= data_out_4[975:960]; end
   9'd445: begin S2_data_out_reg <= data_out_4[991:976]; end
   9'd446: begin S2_data_out_reg <= data_out_4[1007:992]; end
   9'd447: begin S2_data_out_reg <= data_out_4[1023:1008]; end
   9'd448: begin S2_data_out_reg <= data_out_4[1039:1024]; end
   9'd449: begin S2_data_out_reg <= data_out_4[1055:1040]; end
   9'd450: begin S2_data_out_reg <= data_out_4[1071:1056]; end
   9'd451: begin S2_data_out_reg <= data_out_4[1087:1072]; end
   9'd452: begin S2_data_out_reg <= data_out_4[1103:1088]; end
   9'd453: begin S2_data_out_reg <= data_out_4[1119:1104]; end
   9'd454: begin S2_data_out_reg <= data_out_4[1135:1120]; end
   9'd455: begin S2_data_out_reg <= data_out_4[1151:1136]; end
   9'd456: begin S2_data_out_reg <= data_out_4[1167:1152]; end
   9'd457: begin S2_data_out_reg <= data_out_4[1183:1168]; end
   9'd458: begin S2_data_out_reg <= data_out_4[1199:1184]; end
   9'd459: begin S2_data_out_reg <= data_out_4[1215:1200]; end
   9'd460: begin S2_data_out_reg <= data_out_4[1231:1216]; end
   9'd461: begin S2_data_out_reg <= data_out_4[1247:1232]; end
   9'd462: begin S2_data_out_reg <= data_out_4[1263:1248]; end
   9'd463: begin S2_data_out_reg <= data_out_4[1279:1264]; end
   9'd464: begin S2_data_out_reg <= data_out_4[1295:1280]; end
   9'd465: begin S2_data_out_reg <= data_out_4[1311:1296]; end
   9'd466: begin S2_data_out_reg <= data_out_4[1327:1312]; end
   9'd467: begin S2_data_out_reg <= data_out_4[1343:1328]; end
   9'd468: begin S2_data_out_reg <= data_out_4[1359:1344]; end
   9'd469: begin S2_data_out_reg <= data_out_4[1375:1360]; end
   9'd470: begin S2_data_out_reg <= data_out_4[1391:1376]; end
   9'd471: begin S2_data_out_reg <= data_out_4[1407:1392]; end
   9'd472: begin S2_data_out_reg <= data_out_4[1423:1408]; end
   9'd473: begin S2_data_out_reg <= data_out_4[1439:1424]; end
   9'd474: begin S2_data_out_reg <= data_out_4[1455:1440]; end
   9'd475: begin S2_data_out_reg <= data_out_4[1471:1456]; end
   9'd476: begin S2_data_out_reg <= data_out_4[1487:1472]; end
   9'd477: begin S2_data_out_reg <= data_out_4[1503:1488]; end
   9'd478: begin S2_data_out_reg <= data_out_4[1519:1504]; end
   9'd479: begin S2_data_out_reg <= data_out_4[1535:1520]; end
   9'd480: begin S2_data_out_reg <= data_out_4[1551:1536]; end
   9'd481: begin S2_data_out_reg <= data_out_4[1567:1552]; end
   9'd482: begin S2_data_out_reg <= data_out_4[1583:1568]; end
   9'd483: begin S2_data_out_reg <= data_out_4[1599:1584]; end
   9'd484: begin S2_data_out_reg <= data_out_4[1615:1600]; end
   9'd485: begin S2_data_out_reg <= data_out_4[1631:1616]; end
   9'd486: begin S2_data_out_reg <= data_out_4[1647:1632]; end
   9'd487: begin S2_data_out_reg <= data_out_4[1663:1648]; end
   9'd488: begin S2_data_out_reg <= data_out_4[1679:1664]; end
   9'd489: begin S2_data_out_reg <= data_out_4[1695:1680]; end
   9'd490: begin S2_data_out_reg <= data_out_4[1711:1696]; end
   9'd491: begin S2_data_out_reg <= data_out_4[1727:1712]; end
   9'd492: begin S2_data_out_reg <= data_out_4[1743:1728]; end
   9'd493: begin S2_data_out_reg <= data_out_4[1759:1744]; end
   9'd494: begin S2_data_out_reg <= data_out_4[1775:1760]; end
   9'd495: begin S2_data_out_reg <= data_out_4[1791:1776]; end
   9'd496: begin S2_data_out_reg <= data_out_4[1807:1792]; end
   9'd497: begin S2_data_out_reg <= data_out_4[1823:1808]; end
   9'd498: begin S2_data_out_reg <= data_out_4[1839:1824]; end
   9'd499: begin S2_data_out_reg <= data_out_4[1855:1840]; end
   9'd500: begin S2_data_out_reg <= data_out_4[1871:1856]; end
   9'd501: begin S2_data_out_reg <= data_out_4[1887:1872]; end
   9'd502: begin S2_data_out_reg <= data_out_4[1903:1888]; end
   9'd503: begin S2_data_out_reg <= data_out_4[1919:1904]; end
   9'd504: begin S2_data_out_reg <= data_out_4[1935:1920]; end
   9'd505: begin S2_data_out_reg <= data_out_4[1951:1936]; end
   9'd506: begin S2_data_out_reg <= data_out_4[1967:1952]; end
   9'd507: begin S2_data_out_reg <= data_out_4[1983:1968]; end
   9'd508: begin S2_data_out_reg <= data_out_4[1999:1984]; end
   9'd509: begin S2_data_out_reg <= data_out_4[2015:2000]; end
   9'd510: begin S2_data_out_reg <= data_out_4[2031:2016]; end
   9'd511: begin S2_data_out_reg <= data_out_4[2047:2032]; end
       default: begin S2_data_out_reg <= 9'b0; end
   endcase   
end


assign Number_w = Number ;

endmodule