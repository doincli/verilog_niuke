module axi_slave_module#
	(
        /*
C_S_AXI_DATA_WIDTH 表示数据总线的位宽
C_S_AXI_ADDR_WIDTH 表示数据地址的位宽
C_S_AXI_DATA_WIDTH表示数据总线的位宽
C_S_AXI_ADDR_WIDTH表示数据地址的位宽
S_AXI_ACLK ：表示总线时钟
S_AXI_ARESETN：系统复位信号，低电平有效
S_AXI_AWADDR：写地址
S_AXI_AWPROT: 表明传输中数据和命令传输的安全级别和权限
S_AXI_AWVALID：表明写地址和控制数据是否有效
S_AXI_AWREADY：指示从设备准备好接收数据和控制信号
S_AXI_WDATA：写数据
S_AXI_WSTRB:写选通用于指示哪些字节通道传输有效数据几个字节对应几个选通信号bit
S_AXI_WVALID:写有效，该信号写数据和写选通信号是有效的
S_AXI_WREADY:写准备，该信号用于表示从机已经准备好，可以接受写入数据
S_AXI_BRESP:主机接口中的写入响应通道端口
S_AXI_BVALID: 写入响应有效，用来指示写入响应通道正在传输有效数据
S_AXI_BREADY: 响应准备，用于表示主机已经准备好接收写入响应信号
S_AXI_ARADDR: 主机接口读地址通道端口,由主机确定并发起读地址
S_AXI_ARPROT:无论是传输数据还是传输指令都将使用该管脚表明传输的权限和安全级别。
S_AXI_ARVALID: 读地址有效，该信号用于表明通道正在发送有些的读地址数据和控制信息
 S_AXI_ARREADY： 读地址准备，该信号表明从机设备已经准备好，可以接收地址和相关控制信号
S_AXI_RDATA：主机接口读数据通道端口
S_AXI_RRESP：   读取响应，该信号用于指示读取操作的状态
S_AXI_RVALID： 读有效，该信号用于指示通道上正在传输需要的数据
S_AXI_RREADY： 读取准备，该信号用来表示主机已经准备好接收从机响应的读取数据

        */
		parameter                C_S_AXI_ID_WIDTH	    = 1,
		parameter                C_S_AXI_DATA_WIDTH	    = 32,
		parameter                C_S_AXI_ADDR_WIDTH	    = 6,
		parameter                C_S_AXI_AWUSER_WIDTH	= 1,//自定义
		parameter                C_S_AXI_ARUSER_WIDTH	= 1,
        parameter                C_S_AXI_WUSER_WIDTH	= 1,
        parameter                C_S_AXI_RUSER_WIDTH	= 1,
        parameter                C_S_AXI_BUSER_WIDTH	= 1
	)
	(
		input wire                                  S_AXI_ACLK      ,
		input wire                                  S_AXI_ARESETN   ,

		input wire [C_S_AXI_ID_WIDTH-1 : 0]         S_AXI_AWID      ,
		input wire [C_S_AXI_ADDR_WIDTH-1 : 0]       S_AXI_AWADDR    ,
		input wire [7 : 0]                          S_AXI_AWLEN     ,
		input wire [2 : 0]                          S_AXI_AWSIZE    ,
		input wire [1 : 0]                          S_AXI_AWBURST   ,
		input wire                                  S_AXI_AWLOCK    ,
		input wire [3 : 0]                          S_AXI_AWCACHE   ,
		input wire [2 : 0]                          S_AXI_AWPROT    ,
		input wire [3 : 0]                          S_AXI_AWQOS     ,
		input wire [3 : 0]                          S_AXI_AWREGION  ,
		input wire [C_S_AXI_AWUSER_WIDTH-1 : 0]     S_AXI_AWUSER    ,
		input wire                                  S_AXI_AWVALID   ,
		output wire                                 S_AXI_AWREADY   ,

		input wire [C_S_AXI_DATA_WIDTH-1 : 0]       S_AXI_WDATA     ,
		input wire [(C_S_AXI_DATA_WIDTH/8)-1 : 0]   S_AXI_WSTRB     ,
		input wire                                  S_AXI_WLAST     ,
		input wire [C_S_AXI_WUSER_WIDTH-1 : 0]      S_AXI_WUSER     ,
		input wire                                  S_AXI_WVALID    ,
		output wire                                 S_AXI_WREADY    ,

		output wire [C_S_AXI_ID_WIDTH-1 : 0]        S_AXI_BID       ,
		output wire [1 : 0]                         S_AXI_BRESP     ,
		output wire [C_S_AXI_BUSER_WIDTH-1 : 0]     S_AXI_BUSER     ,
		output wire                                 S_AXI_BVALID    ,
		input wire                                  S_AXI_BREADY    ,

		input wire [C_S_AXI_ID_WIDTH-1 : 0]         S_AXI_ARID      ,
		input wire [C_S_AXI_ADDR_WIDTH-1 : 0]       S_AXI_ARADDR    ,
		input wire [7 : 0]                          S_AXI_ARLEN     ,
		input wire [2 : 0]                          S_AXI_ARSIZE    ,
		input wire [1 : 0]                          S_AXI_ARBURST   ,
		input wire                                  S_AXI_ARLOCK    ,
		input wire [3 : 0]                          S_AXI_ARCACHE   ,
		input wire [2 : 0]                          S_AXI_ARPROT    ,
		input wire [3 : 0]                          S_AXI_ARQOS     ,
		input wire [3 : 0]                          S_AXI_ARREGION  ,
		input wire [C_S_AXI_ARUSER_WIDTH-1 : 0]     S_AXI_ARUSER    ,
		input wire                                  S_AXI_ARVALID   ,
		output wire                                 S_AXI_ARREADY   ,

		output wire [C_S_AXI_ID_WIDTH-1 : 0]        S_AXI_RID       ,
		output wire [C_S_AXI_DATA_WIDTH-1 : 0]      S_AXI_RDATA     ,
		output wire [1 : 0]                         S_AXI_RRESP     ,
		output wire                                 S_AXI_RLAST     ,
		output wire [C_S_AXI_RUSER_WIDTH-1 : 0]     S_AXI_RUSER     ,
		output wire                                 S_AXI_RVALID    ,
		input wire                                  S_AXI_RREADY    
);

/**********************参数***************************/

/**********************状态机*************************/

/**********************寄存器*************************/
reg [C_S_AXI_ADDR_WIDTH-1 : 0]  r_awaddr                                ;
reg [7 : 0]                     r_awlen                                 ;
reg                             r_awready                               ;
reg                             r_wready                                ;
reg                             r_arready                               ;
reg [C_S_AXI_ADDR_WIDTH-1 : 0]  r_araddr                                ;
reg [7 : 0]                     r_arlen                                 ;
reg [7 : 0]                     r_read_cnt                              ;
reg                             r_rvalid                                ;
reg                             r_rvalid_1b                             ;
reg                             r_rvalid_2b                             ;
reg                             r_bvalid                                ;

reg [C_S_AXI_DATA_WIDTH-1 : 0]  r_ram[0 : 255]                          ;
reg [7:0]                       r_ram_addr                              ;
reg [7:0]                       r_ram_addr_1b                           ;   
reg [C_S_AXI_DATA_WIDTH-1 : 0]  r_ram_write_data                        ;
reg [C_S_AXI_DATA_WIDTH-1 : 0]  r_ram_read_data                         ;
reg                             r_ram_rh_wl                             ;
reg                             r_ram_en                                ;

/**********************网表型*************************/ 
wire                w_aw_active                                         ;
wire                w_w_active                                          ;
wire                w_b_active                                          ;
wire                w_ar_active                                         ;
wire                w_r_active                                          ;
wire                w_rst                                               ;

/**********************组合逻辑***********************/
assign              w_aw_active     = S_AXI_AWVALID   & S_AXI_AWREADY   ;
assign              w_w_active      = S_AXI_WVALID    & S_AXI_WREADY    ;
assign              w_b_active      = S_AXI_BVALID    & S_AXI_BREADY    ;
assign              w_ar_active     = S_AXI_ARVALID   & S_AXI_ARREADY   ;
assign              w_r_active      = S_AXI_RVALID    & S_AXI_RREADY    ;
assign              S_AXI_AWREADY   = r_awready                         ;
assign              S_AXI_WREADY    = r_wready                          ;
assign              S_AXI_ARREADY   = r_arready                         ;
assign              w_rst           = ~S_AXI_ARESETN                    ;

assign              S_AXI_RID       = 'd0                               ;
assign              S_AXI_RDATA     = r_ram_read_data                   ;
assign              S_AXI_RRESP     = 'd0                               ;
assign              S_AXI_RLAST     = (r_read_cnt == r_arlen - 1) ? 
                                      w_r_active : 1'b0                 ; 
assign              S_AXI_RUSER     = 'd0                               ;
assign              S_AXI_RVALID    = r_rvalid_2b                       ;
assign              S_AXI_BID       = 'd0                               ;
assign              S_AXI_BRESP     = 'd0                               ;
assign              S_AXI_BUSER     = 'd0                               ;
assign              S_AXI_BVALID    = r_bvalid                          ;
/**********************例化***************************/

/**********************进程***************************/
//写地址
always@(posedge S_AXI_ACLK)
    if(w_aw_active)
        r_awaddr <= S_AXI_AWADDR;
    else 
        r_awaddr <= r_awaddr;

//写长度
always@(posedge S_AXI_ACLK)
    if(w_aw_active)
        r_awlen <= S_AXI_AWLEN;
    // else if()
    else 
        r_awlen <= r_awlen;

//写地址准备信号
always@(posedge S_AXI_ACLK)
    if(w_rst || S_AXI_WLAST)
        r_awready <= 'd1;
    else if(w_aw_active)   
        r_awready <= 'd0;
    else    
        r_awready <= r_awready;

//写数据准备信号
always@(posedge S_AXI_ACLK)
    if(w_aw_active)
        r_wready <= 'd1;
    else if(S_AXI_WLAST)
        r_wready <= 'd0;
    else 
        r_wready <= r_wready;

//ram核心写
always@(posedge S_AXI_ACLK)
    if(!r_ram_rh_wl) 
        r_ram[r_ram_addr_1b] <= r_ram_en ? r_ram_write_data : r_ram[r_ram_addr];
    else 
        r_ram[r_ram_addr_1b] <= r_ram[r_ram_addr_1b];

//ram核心读
always@(posedge S_AXI_ACLK)
    if(r_ram_rh_wl)
        r_ram_read_data <= r_ram[r_ram_addr_1b] ;  
    else 
        r_ram_read_data <= r_ram_read_data   ;

//ram地址
always@(posedge S_AXI_ACLK)
    if(w_rst || S_AXI_WLAST || S_AXI_RLAST)
        r_ram_addr <= 'd0;
    else if(w_aw_active)
        r_ram_addr <= S_AXI_AWADDR[7:0];
    else if(w_ar_active)
        r_ram_addr <= S_AXI_ARADDR[7:0];
    else if(w_w_active || (r_rvalid & S_AXI_RREADY))
        r_ram_addr <= r_ram_addr + 1;
    else 
        r_ram_addr <= r_ram_addr;

//ram地址打一拍
always@(posedge S_AXI_ACLK)
    r_ram_addr_1b <= r_ram_addr;

//ram写端口
always@(posedge S_AXI_ACLK)
    if(w_w_active)
        r_ram_write_data <= S_AXI_WDATA         ;
    else    
        r_ram_write_data <= r_ram_write_data    ;

//ram读写控制
always@(posedge S_AXI_ACLK)
    if(w_ar_active)
        r_ram_rh_wl <= 'd1;
    else if(w_aw_active)
        r_ram_rh_wl <= 'd0;
    else 
        r_ram_rh_wl <= r_ram_rh_wl;

//ram写使能
always@(posedge S_AXI_ACLK)
    if(w_w_active)
        r_ram_en <= 'd1;
    else
        r_ram_en <= 'd0;



always@(posedge S_AXI_ACLK)
    if(w_rst || S_AXI_RLAST)
        r_arready <= 'd1;
    else if(w_ar_active)
        r_arready <= 'd0;
    else 
        r_arready <= r_arready;

 
always@(posedge S_AXI_ACLK)
    if(w_ar_active)
        r_araddr <= S_AXI_ARADDR;
    else 
        r_araddr <= r_araddr;

always@(posedge S_AXI_ACLK)
    if(w_ar_active)
        r_arlen <= S_AXI_ARLEN; 
    else 
        r_arlen <= r_arlen;

always@(posedge S_AXI_ACLK)
    if(w_rst || S_AXI_RLAST)
        r_read_cnt <= 'd0;
    else if(w_r_active)
        r_read_cnt <= r_read_cnt + 1;
    else 
        r_read_cnt <= r_read_cnt;

always@(posedge S_AXI_ACLK)
    if(w_rst || S_AXI_RLAST)
        r_rvalid <= 'd0;
    else if(w_ar_active)
        r_rvalid <= 'd1;
    else 
        r_rvalid <= r_rvalid;

always@(posedge S_AXI_ACLK)
    if(S_AXI_RLAST)
        r_rvalid_1b <= 'd0;
    else 
        r_rvalid_1b <= r_rvalid;

always@(posedge S_AXI_ACLK)
    if(S_AXI_RLAST)
        r_rvalid_2b <= 'd0;
    else 
        r_rvalid_2b <= r_rvalid_1b;

always@(posedge S_AXI_ACLK)
    if(S_AXI_WLAST)
        r_bvalid <= 'd1;
    else if(w_b_active)
        r_bvalid <= 'd0;
    else 
        r_bvalid <= r_bvalid;
endmodule
